module pipeline_regs (
    input logic clk,
    input logic reset
);
    // Pipeline registers will be added in later milestones
endmodule
